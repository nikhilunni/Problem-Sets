// Design a circuit that divides a 4-bit signed binary number (in)
// by 3 to produce a 3-bit signed binary number (out).  Note that
// integer division rounds toward zero for both positive and negative
// numbers (e.g., -5/3 is -1).

module sdiv3(out, in);
   output [2:0] out;
   input  [3:0]	in;
   
endmodule // sdiv3

